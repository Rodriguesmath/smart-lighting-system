module maquina_principal (
    input logic clk, rst, a, b, c, d,
    output logic led, saida
);

  // Implementação da máquina de estados principal
  // ...

endmodule