module module_2 #(
    parameter AUTO_SHUTDOWN_T = 30000
)(
    input wire clk, rst,
    input logic infravermelho,
    output logic C
);

  // Implementação da máquina de estados para o controle do tempo da lâmpada
  // ...

endmodule